magic
tech sky130A
magscale 1 2
timestamp 1671089792
<< nwell >>
rect 1066 87301 38862 87622
rect 1066 86213 38862 86779
rect 1066 85125 38862 85691
rect 1066 84037 38862 84603
rect 1066 82949 38862 83515
rect 1066 81861 38862 82427
rect 1066 80773 38862 81339
rect 1066 79685 38862 80251
rect 1066 78597 38862 79163
rect 1066 77509 38862 78075
rect 1066 76421 38862 76987
rect 1066 75333 38862 75899
rect 1066 74245 38862 74811
rect 1066 73157 38862 73723
rect 1066 72069 38862 72635
rect 1066 70981 38862 71547
rect 1066 69893 38862 70459
rect 1066 68805 38862 69371
rect 1066 67717 38862 68283
rect 1066 66629 38862 67195
rect 1066 65541 38862 66107
rect 1066 64453 38862 65019
rect 1066 63365 38862 63931
rect 1066 62277 38862 62843
rect 1066 61189 38862 61755
rect 1066 60101 38862 60667
rect 1066 59013 38862 59579
rect 1066 57925 38862 58491
rect 1066 56837 38862 57403
rect 1066 55749 38862 56315
rect 1066 54661 38862 55227
rect 1066 53573 38862 54139
rect 1066 52485 38862 53051
rect 1066 51397 38862 51963
rect 1066 50309 38862 50875
rect 1066 49221 38862 49787
rect 1066 48133 38862 48699
rect 1066 47045 38862 47611
rect 1066 45957 38862 46523
rect 1066 44869 38862 45435
rect 1066 43781 38862 44347
rect 1066 42693 38862 43259
rect 1066 41605 38862 42171
rect 1066 40517 38862 41083
rect 1066 39429 38862 39995
rect 1066 38341 38862 38907
rect 1066 37253 38862 37819
rect 1066 36165 38862 36731
rect 1066 35077 38862 35643
rect 1066 33989 38862 34555
rect 1066 32901 38862 33467
rect 1066 31813 38862 32379
rect 1066 30725 38862 31291
rect 1066 29637 38862 30203
rect 1066 28549 38862 29115
rect 1066 27461 38862 28027
rect 1066 26373 38862 26939
rect 1066 25285 38862 25851
rect 1066 24197 38862 24763
rect 1066 23109 38862 23675
rect 1066 22021 38862 22587
rect 1066 20933 38862 21499
rect 1066 19845 38862 20411
rect 1066 18757 38862 19323
rect 1066 17669 38862 18235
rect 1066 16581 38862 17147
rect 1066 15493 38862 16059
rect 1066 14405 38862 14971
rect 1066 13317 38862 13883
rect 1066 12229 38862 12795
rect 1066 11141 38862 11707
rect 1066 10053 38862 10619
rect 1066 8965 38862 9531
rect 1066 7877 38862 8443
rect 1066 6789 38862 7355
rect 1066 5701 38862 6267
rect 1066 4613 38862 5179
rect 1066 3525 38862 4091
rect 1066 2437 38862 3003
<< obsli1 >>
rect 1104 2159 38824 87601
<< obsm1 >>
rect 1104 2128 38824 87712
<< metal2 >>
rect 1214 89200 1270 90000
rect 2778 89200 2834 90000
rect 4342 89200 4398 90000
rect 5906 89200 5962 90000
rect 7470 89200 7526 90000
rect 9034 89200 9090 90000
rect 10598 89200 10654 90000
rect 12162 89200 12218 90000
rect 13726 89200 13782 90000
rect 15290 89200 15346 90000
rect 16854 89200 16910 90000
rect 18418 89200 18474 90000
rect 19982 89200 20038 90000
rect 21546 89200 21602 90000
rect 23110 89200 23166 90000
rect 24674 89200 24730 90000
rect 26238 89200 26294 90000
rect 27802 89200 27858 90000
rect 29366 89200 29422 90000
rect 30930 89200 30986 90000
rect 32494 89200 32550 90000
rect 34058 89200 34114 90000
rect 35622 89200 35678 90000
rect 37186 89200 37242 90000
rect 38750 89200 38806 90000
rect 9954 0 10010 800
rect 29918 0 29974 800
<< obsm2 >>
rect 1326 89144 2722 89298
rect 2890 89144 4286 89298
rect 4454 89144 5850 89298
rect 6018 89144 7414 89298
rect 7582 89144 8978 89298
rect 9146 89144 10542 89298
rect 10710 89144 12106 89298
rect 12274 89144 13670 89298
rect 13838 89144 15234 89298
rect 15402 89144 16798 89298
rect 16966 89144 18362 89298
rect 18530 89144 19926 89298
rect 20094 89144 21490 89298
rect 21658 89144 23054 89298
rect 23222 89144 24618 89298
rect 24786 89144 26182 89298
rect 26350 89144 27746 89298
rect 27914 89144 29310 89298
rect 29478 89144 30874 89298
rect 31042 89144 32438 89298
rect 32606 89144 34002 89298
rect 34170 89144 35566 89298
rect 35734 89144 37130 89298
rect 37298 89144 38694 89298
rect 1270 856 38804 89144
rect 1270 800 9898 856
rect 10066 800 29862 856
rect 30030 800 38804 856
<< obsm3 >>
rect 4210 2143 35246 87617
<< metal4 >>
rect 4208 2128 4528 87632
rect 19568 2128 19888 87632
rect 34928 2128 35248 87632
<< obsm4 >>
rect 11835 6835 12637 72045
<< labels >>
rlabel metal2 s 9954 0 10010 800 6 clock
port 1 nsew signal input
rlabel metal2 s 1214 89200 1270 90000 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 26238 89200 26294 90000 6 io_in[10]
port 3 nsew signal input
rlabel metal2 s 27802 89200 27858 90000 6 io_in[11]
port 4 nsew signal input
rlabel metal2 s 29366 89200 29422 90000 6 io_in[12]
port 5 nsew signal input
rlabel metal2 s 30930 89200 30986 90000 6 io_in[13]
port 6 nsew signal input
rlabel metal2 s 32494 89200 32550 90000 6 io_in[14]
port 7 nsew signal input
rlabel metal2 s 34058 89200 34114 90000 6 io_in[15]
port 8 nsew signal input
rlabel metal2 s 35622 89200 35678 90000 6 io_in[16]
port 9 nsew signal input
rlabel metal2 s 37186 89200 37242 90000 6 io_in[17]
port 10 nsew signal input
rlabel metal2 s 38750 89200 38806 90000 6 io_in[18]
port 11 nsew signal input
rlabel metal2 s 5906 89200 5962 90000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 10598 89200 10654 90000 6 io_in[2]
port 13 nsew signal input
rlabel metal2 s 15290 89200 15346 90000 6 io_in[3]
port 14 nsew signal input
rlabel metal2 s 16854 89200 16910 90000 6 io_in[4]
port 15 nsew signal input
rlabel metal2 s 18418 89200 18474 90000 6 io_in[5]
port 16 nsew signal input
rlabel metal2 s 19982 89200 20038 90000 6 io_in[6]
port 17 nsew signal input
rlabel metal2 s 21546 89200 21602 90000 6 io_in[7]
port 18 nsew signal input
rlabel metal2 s 23110 89200 23166 90000 6 io_in[8]
port 19 nsew signal input
rlabel metal2 s 24674 89200 24730 90000 6 io_in[9]
port 20 nsew signal input
rlabel metal2 s 2778 89200 2834 90000 6 io_oeb[0]
port 21 nsew signal output
rlabel metal2 s 7470 89200 7526 90000 6 io_oeb[1]
port 22 nsew signal output
rlabel metal2 s 12162 89200 12218 90000 6 io_oeb[2]
port 23 nsew signal output
rlabel metal2 s 4342 89200 4398 90000 6 io_out[0]
port 24 nsew signal output
rlabel metal2 s 9034 89200 9090 90000 6 io_out[1]
port 25 nsew signal output
rlabel metal2 s 13726 89200 13782 90000 6 io_out[2]
port 26 nsew signal output
rlabel metal2 s 29918 0 29974 800 6 reset
port 27 nsew signal input
rlabel metal4 s 4208 2128 4528 87632 6 vccd1
port 28 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 87632 6 vccd1
port 28 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 87632 6 vssd1
port 29 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 90000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1694362
string GDS_FILE /home/abdulkadr/Desktop/caravel_first/openlane/oto_pilot/runs/22_12_15_10_35/results/signoff/oto_pilot.magic.gds
string GDS_START 376474
<< end >>

