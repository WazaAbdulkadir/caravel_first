VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO oto_pilot
  CLASS BLOCK ;
  FOREIGN oto_pilot ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 450.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END clock
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 446.000 6.350 450.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 446.000 131.470 450.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 446.000 139.290 450.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 446.000 147.110 450.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 446.000 154.930 450.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 446.000 162.750 450.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 446.000 170.570 450.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 446.000 178.390 450.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 446.000 186.210 450.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 446.000 194.030 450.000 ;
    END
  END io_in[18]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 446.000 29.810 450.000 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 446.000 53.270 450.000 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 446.000 76.730 450.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 446.000 84.550 450.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 446.000 92.370 450.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 446.000 100.190 450.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 446.000 108.010 450.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 446.000 115.830 450.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 446.000 123.650 450.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 446.000 14.170 450.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 446.000 37.630 450.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 446.000 61.090 450.000 ;
    END
  END io_oeb[2]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 446.000 21.990 450.000 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 446.000 45.450 450.000 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 446.000 68.910 450.000 ;
    END
  END io_out[2]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 438.160 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 438.160 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 436.505 194.310 438.110 ;
        RECT 5.330 431.065 194.310 433.895 ;
        RECT 5.330 425.625 194.310 428.455 ;
        RECT 5.330 420.185 194.310 423.015 ;
        RECT 5.330 414.745 194.310 417.575 ;
        RECT 5.330 409.305 194.310 412.135 ;
        RECT 5.330 403.865 194.310 406.695 ;
        RECT 5.330 398.425 194.310 401.255 ;
        RECT 5.330 392.985 194.310 395.815 ;
        RECT 5.330 387.545 194.310 390.375 ;
        RECT 5.330 382.105 194.310 384.935 ;
        RECT 5.330 376.665 194.310 379.495 ;
        RECT 5.330 371.225 194.310 374.055 ;
        RECT 5.330 365.785 194.310 368.615 ;
        RECT 5.330 360.345 194.310 363.175 ;
        RECT 5.330 354.905 194.310 357.735 ;
        RECT 5.330 349.465 194.310 352.295 ;
        RECT 5.330 344.025 194.310 346.855 ;
        RECT 5.330 338.585 194.310 341.415 ;
        RECT 5.330 333.145 194.310 335.975 ;
        RECT 5.330 327.705 194.310 330.535 ;
        RECT 5.330 322.265 194.310 325.095 ;
        RECT 5.330 316.825 194.310 319.655 ;
        RECT 5.330 311.385 194.310 314.215 ;
        RECT 5.330 305.945 194.310 308.775 ;
        RECT 5.330 300.505 194.310 303.335 ;
        RECT 5.330 295.065 194.310 297.895 ;
        RECT 5.330 289.625 194.310 292.455 ;
        RECT 5.330 284.185 194.310 287.015 ;
        RECT 5.330 278.745 194.310 281.575 ;
        RECT 5.330 273.305 194.310 276.135 ;
        RECT 5.330 267.865 194.310 270.695 ;
        RECT 5.330 262.425 194.310 265.255 ;
        RECT 5.330 256.985 194.310 259.815 ;
        RECT 5.330 251.545 194.310 254.375 ;
        RECT 5.330 246.105 194.310 248.935 ;
        RECT 5.330 240.665 194.310 243.495 ;
        RECT 5.330 235.225 194.310 238.055 ;
        RECT 5.330 229.785 194.310 232.615 ;
        RECT 5.330 224.345 194.310 227.175 ;
        RECT 5.330 218.905 194.310 221.735 ;
        RECT 5.330 213.465 194.310 216.295 ;
        RECT 5.330 208.025 194.310 210.855 ;
        RECT 5.330 202.585 194.310 205.415 ;
        RECT 5.330 197.145 194.310 199.975 ;
        RECT 5.330 191.705 194.310 194.535 ;
        RECT 5.330 186.265 194.310 189.095 ;
        RECT 5.330 180.825 194.310 183.655 ;
        RECT 5.330 175.385 194.310 178.215 ;
        RECT 5.330 169.945 194.310 172.775 ;
        RECT 5.330 164.505 194.310 167.335 ;
        RECT 5.330 159.065 194.310 161.895 ;
        RECT 5.330 153.625 194.310 156.455 ;
        RECT 5.330 148.185 194.310 151.015 ;
        RECT 5.330 142.745 194.310 145.575 ;
        RECT 5.330 137.305 194.310 140.135 ;
        RECT 5.330 131.865 194.310 134.695 ;
        RECT 5.330 126.425 194.310 129.255 ;
        RECT 5.330 120.985 194.310 123.815 ;
        RECT 5.330 115.545 194.310 118.375 ;
        RECT 5.330 110.105 194.310 112.935 ;
        RECT 5.330 104.665 194.310 107.495 ;
        RECT 5.330 99.225 194.310 102.055 ;
        RECT 5.330 93.785 194.310 96.615 ;
        RECT 5.330 88.345 194.310 91.175 ;
        RECT 5.330 82.905 194.310 85.735 ;
        RECT 5.330 77.465 194.310 80.295 ;
        RECT 5.330 72.025 194.310 74.855 ;
        RECT 5.330 66.585 194.310 69.415 ;
        RECT 5.330 61.145 194.310 63.975 ;
        RECT 5.330 55.705 194.310 58.535 ;
        RECT 5.330 50.265 194.310 53.095 ;
        RECT 5.330 44.825 194.310 47.655 ;
        RECT 5.330 39.385 194.310 42.215 ;
        RECT 5.330 33.945 194.310 36.775 ;
        RECT 5.330 28.505 194.310 31.335 ;
        RECT 5.330 23.065 194.310 25.895 ;
        RECT 5.330 17.625 194.310 20.455 ;
        RECT 5.330 12.185 194.310 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 194.120 438.005 ;
      LAYER met1 ;
        RECT 5.520 10.640 194.120 438.560 ;
      LAYER met2 ;
        RECT 6.630 445.720 13.610 446.490 ;
        RECT 14.450 445.720 21.430 446.490 ;
        RECT 22.270 445.720 29.250 446.490 ;
        RECT 30.090 445.720 37.070 446.490 ;
        RECT 37.910 445.720 44.890 446.490 ;
        RECT 45.730 445.720 52.710 446.490 ;
        RECT 53.550 445.720 60.530 446.490 ;
        RECT 61.370 445.720 68.350 446.490 ;
        RECT 69.190 445.720 76.170 446.490 ;
        RECT 77.010 445.720 83.990 446.490 ;
        RECT 84.830 445.720 91.810 446.490 ;
        RECT 92.650 445.720 99.630 446.490 ;
        RECT 100.470 445.720 107.450 446.490 ;
        RECT 108.290 445.720 115.270 446.490 ;
        RECT 116.110 445.720 123.090 446.490 ;
        RECT 123.930 445.720 130.910 446.490 ;
        RECT 131.750 445.720 138.730 446.490 ;
        RECT 139.570 445.720 146.550 446.490 ;
        RECT 147.390 445.720 154.370 446.490 ;
        RECT 155.210 445.720 162.190 446.490 ;
        RECT 163.030 445.720 170.010 446.490 ;
        RECT 170.850 445.720 177.830 446.490 ;
        RECT 178.670 445.720 185.650 446.490 ;
        RECT 186.490 445.720 193.470 446.490 ;
        RECT 6.350 4.280 194.020 445.720 ;
        RECT 6.350 4.000 49.490 4.280 ;
        RECT 50.330 4.000 149.310 4.280 ;
        RECT 150.150 4.000 194.020 4.280 ;
      LAYER met3 ;
        RECT 21.050 10.715 176.230 438.085 ;
      LAYER met4 ;
        RECT 59.175 34.175 63.185 360.225 ;
  END
END oto_pilot
END LIBRARY

